module not_gate( Out, In );
    input In;
    output Out;

    assign Out = ~In;
endmodule
